`include "lnrv_def.v"
module  lnrv_idu_decode
(
    // 指令输入
    input[31 : 0]                       ir,

    output[4 : 0]                       dec_rs1_idx,
    output[4 : 0]                       dec_rs2_idx,
    output[4 : 0]                       dec_rd_idx,
    output[11 : 0]                      dec_csr_idx,
    output[31 : 0]                      dec_imm,

    // 指令长度指示
    output                              dec_rv32,
    output                              dec_rv16,

    input                               d_mode,

    // 非法指令
    output                              dec_ilegl_instr,

    output[`DEC_OP_BUS_WIDTH - 1 : 0]   dec_op_bus,
    output                              dec_rglr_instr,     // 常规指令
    output                              dec_lsu_instr,      // load and store指令
    output                              dec_csr_instr,
    output                              dec_brch_instr,     // 分支相关指令
    output                              dec_mdv_instr,      // 乘除法相关指令
    output                              dec_sys_instr,      // 系统相关指令
    output                              dec_amo_instr,
    output                              dec_fpu_instr
);


wire[6 : 0]                         opcode;
wire                                opcode_is_0110111;
wire                                opcode_is_0010111;
wire                                opcode_is_1101111;
wire                                opcode_is_1100111;
wire                                opcode_is_1100011;
wire                                opcode_is_0000011;
wire                                opcode_is_0100011;
wire                                opcode_is_0010011;
wire                                opcode_is_0110011;
wire                                opcode_is_0001111;
wire                                opcode_is_1110011;
wire                                opcode_is_0101111;
wire                                funct7_is_0001000;


wire[2 : 0]                         funct3;
wire	                            funct3_is_000;
wire	                            funct3_is_001;
wire	                            funct3_is_010;
wire	                            funct3_is_011;
wire	                            funct3_is_100;
wire	                            funct3_is_101;
wire	                            funct3_is_110;
wire	                            funct3_is_111;

wire[6 : 0]                         funct7;
wire	                            funct7_is_0000000;
wire	                            funct7_is_0100000;
wire	                            funct7_is_0000001;

// 指令类型
wire                                instr_is_u_type;
wire                                instr_is_i_type;
wire                                instr_is_s_type;
wire                                instr_is_b_type;
wire                                instr_is_j_type;
wire                                instr_is_r_type;

// 具体指令
// 常规指令
wire                                instr_is_add;
wire                                instr_is_addi;
wire                                instr_is_and;
wire                                instr_is_andi;
wire                                instr_is_auipc;
wire                                instr_is_or;
wire                                instr_is_ori;
wire                                instr_is_xor;
wire                                instr_is_xori;
wire                                instr_is_sll;
wire                                instr_is_slli;
wire                                instr_is_slt;
wire                                instr_is_slti;
wire                                instr_is_sltiu;
wire                                instr_is_sltu;
wire                                instr_is_sra;
wire                                instr_is_srai;
wire                                instr_is_srl;
wire                                instr_is_srli;
wire                                instr_is_sub;
wire                                instr_is_lui;

// csr相关指令
wire                                instr_is_csrrc;
wire                                instr_is_csrrci;
wire                                instr_is_csrrw;
wire                                instr_is_csrrwi;
wire                                instr_is_csrrs;
wire                                instr_is_csrrsi;

// 分支相关指令
wire                                instr_is_beq;
wire                                instr_is_bge;
wire                                instr_is_bgeu;
wire                                instr_is_blt;
wire                                instr_is_bltu;
wire                                instr_is_bne;
wire                                instr_is_jal;
wire                                instr_is_jalr;

// 系统相关指令
wire                                instr_is_ebreak;
wire                                instr_is_ecall;
wire                                instr_is_dret;
wire                                instr_is_mret;
wire                                instr_is_fence;
wire                                instr_is_fencei;
wire                                instr_is_wfi;

// load and store相关指令
wire                                instr_is_lb;
wire                                instr_is_lbu;
wire                                instr_is_lh;
wire                                instr_is_lhu;
wire                                instr_is_lrw;
wire                                instr_is_lw;
wire                                instr_is_scw;
wire                                instr_is_sb;
wire                                instr_is_sh;
wire                                instr_is_sw;

wire                                instr_is_div;
wire                                instr_is_divu;
wire                                instr_is_mul;
wire                                instr_is_mulh;
wire                                instr_is_mulhsu;
wire                                instr_is_mulhu;
wire                                instr_is_rem;
wire                                instr_is_remu;



// 不同类型指令的立即数位置不同
wire[31 : 0]                        i_type_imm;
wire[31 : 0]                        i_type_shamt;
wire[31 : 0]                        i_type_zimm;
wire[31 : 0]                        b_type_bxx_imm;
wire[31 : 0]                        b_type_jal_imm;
wire[31 : 0]                        s_type_imm;
wire[31 : 0]                        u_type_imm;
wire[31 : 0]                        j_type_imm;

wire                                sel_i_type_imm;
wire                                sel_i_type_shamt;
wire                                sel_i_type_zimm;
wire                                sel_b_type_bxx_imm;
wire                                sel_b_type_jal_imm;
wire                                sel_s_type_imm;
wire                                sel_u_type_imm;


wire[4 : 0]                         rs1_idx;
wire[4 : 0]                         rs2_idx;
wire[4 : 0]                         rd_idx;
wire[11 : 0]                        csr_idx;

wire[`RGLR_OP_BUS_WIDTH - 1 : 0]    rglr_op_bus;
wire[`BRCH_OP_BUS_WIDTH - 1 : 0]    brch_op_bus;
wire[`SYS_OP_BUS_WIDTH - 1 : 0]     sys_op_bus;
wire[`LSU_OP_BUS_WIDTH - 1 : 0]     lsu_op_bus;
wire[`CSR_OP_BUS_WIDTH - 1 : 0]     csr_op_bus;
wire[`MDV_OP_BUS_WIDTH - 1 : 0]     mdv_op_bus;
wire[`DEC_OP_BUS_WIDTH : 0]         dec_op_bus_mux;

wire                                ilegl_dret;
wire                                legl_dret;
wire                                ilegl_shamt;
wire                                ilegl_sxxi;
wire                                legl_exu;
wire                                ilegl_exu;

// 首先从指令中解析opcode、funct3以及funct7，并分类
assign      opcode = `GET_INSTR_OPCODE(ir);
assign      opcode_is_0110111 = (opcode == 7'b0110111);
assign      opcode_is_0010111 = (opcode == 7'b0010111);
assign      opcode_is_1101111 = (opcode == 7'b1101111);
assign      opcode_is_1100111 = (opcode == 7'b1100111);
assign      opcode_is_1100011 = (opcode == 7'b1100011);
assign      opcode_is_0000011 = (opcode == 7'b0000011);
assign      opcode_is_0100011 = (opcode == 7'b0100011);
assign      opcode_is_0010011 = (opcode == 7'b0010011);
assign      opcode_is_0110011 = (opcode == 7'b0110011);
assign      opcode_is_0001111 = (opcode == 7'b0001111);
assign      opcode_is_1110011 = (opcode == 7'b1110011);
assign      opcode_is_0101111 = (opcode == 7'b0101111);


assign      funct3 = `GET_INSTR_FUNCT3(ir);
assign      funct3_is_000 = (funct3 == 3'b000);
assign      funct3_is_001 = (funct3 == 3'b001);
assign      funct3_is_010 = (funct3 == 3'b010);
assign      funct3_is_011 = (funct3 == 3'b011);
assign      funct3_is_100 = (funct3 == 3'b100);
assign      funct3_is_101 = (funct3 == 3'b101);
assign      funct3_is_110 = (funct3 == 3'b110);
assign      funct3_is_111 = (funct3 == 3'b111);

assign      funct7 = `GET_INSTR_FUNCT7(ir);
assign      funct7_is_0000000 = (funct7 == 7'b0000000);
assign      funct7_is_0100000 = (funct7 == 7'b0100000);
assign      funct7_is_0000001 = (funct7 == 7'b0000001);
assign      funct7_is_0001000 = (funct7 == 7'b0001000);


// 判断指令类型
assign      instr_is_u_type =   opcode_is_0110111 | 
                                opcode_is_0010111;

assign      instr_is_j_type =   opcode_is_1101111;

assign      instr_is_i_type =   opcode_is_1100111 | 
                                opcode_is_0000011 | 
                                opcode_is_0010011 | 
                                opcode_is_0001111 | 
                                opcode_is_1110011;

assign      instr_is_b_type =   opcode_is_1100011;
assign      instr_is_s_type =   opcode_is_0100011;
assign      instr_is_r_type =   opcode_is_0110011;

// 提取寄存器索引
assign      rs1_idx = ir[19 : 15];
assign      rs2_idx = ir[24 : 20];
assign      rd_idx  = ir[11 : 7];
assign      csr_idx = ir[31 : 20];

/*
    add 加，R-Type，RV32I and RV64I，		x[rd] = x[rs1] + x[rs2]，忽略算术溢出
    +----------------------------------------------------------------------------+
    |31				 25|24		20|19		15|14	12|11		   7|6			0|
    +------------------+----------+-----------+-------+-------------+------------+
    |		0000000	   |    rs2	  |    rs1    |  000  | 	rd		|   0110011  |
    +----------------------------------------------------------------------------+
*/
assign      instr_is_add = opcode_is_0110011 & funct3_is_000 & funct7_is_0000000;

/*
    addi 加立即数，I-Type，RV32I and RV64I，	x[rd] = x[rs1] + sext[imm[11 : 0]];
    加符号位扩展的立即数加到寄存器x[rs1]上，并将结果写入x[rd]，忽略算术溢出
    +----------------------------------------------------------------------------+
    |31				 			20|19		15|14	12|11		   7|6			0|
    +-----------------------------+-----------+-------+-------------+------------+
    |		imm[11:0]			  |    rs1    |  000  | 	rd		|   0010011  |
    +----------------------------------------------------------------------------+
*/
assign      instr_is_addi = opcode_is_0010011 & funct3_is_000;

/*
	and 与, R-Type, RV32I and RV64I, 					x[rd] = x[rs1] & x[rs2];
	将寄存器x[rs1]和寄存器x[rs2]位与的结果写入x[rd]寄存器.
	+----------------------------------------------------------------------------+
	|31				 25|24		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|		0000000	   |    rs2	  |    rs1    |  111  | 	rd		|   0110011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_and = opcode_is_0110011 & funct3_is_111 & funct7_is_0000000;

/*
    andi 与立即数, I-Type, RV32I and RV64I, x[rd] = x[rs1] & sext(imm[11 : 0]);
    把符号位扩展的立即数和寄存器x[rs1]位与的结果写入x[rd]寄存器.
    +----------------------------------------------------------------------------+
    |31				 			20|19		15|14	12|11		   7|6			0|
    +-----------------------------+-----------+-------+-------------+------------+
    |		imm[11:0]			  |    rs1    |  111  | 	rd		|   0010011  |
    +----------------------------------------------------------------------------+
*/
assign      instr_is_andi = opcode_is_0010011 & funct3_is_111;

/* 
	auipc PC加立即数, U-Type, x[rd] = PC + sext(imm[31 : 12] << 12);
	把符号位扩展的20位(左移12位)立即数加到PC上，并将结果写入x[rd].
	+----------------------------------------------------------------------------+
	|31				 								12|11		   7|6			0|
	+-------------------------------------------------+-------------+------------+
	|					imm[31:12]		  			  | 	rd		|  0010111   |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_auipc = opcode_is_0010111;

/*
    beq	相等时分支, B-Type, RV32I and RV64I, if(x[rs1] == x[rs2])	pc += sext(imm);
    若寄存器x[rs1]和寄存器x[rs2]的值相等，把pc的值设置为当前值加上符号位扩展的立即数;
        ----------------------------------------------------------------------------
    |31              25|24      20|19		15|14	12|11		   7|6			0|
        ------------------ ---------- ----------- ------- ------------- ------------
    |	imm[12|10:5]   |    rs2	  |    rs1    |  000  | imm[4:1|11] |   1100011  |
        ----------------------------------------------------------------------------
*/
assign      instr_is_beq = opcode_is_1100011 & funct3_is_000;

/*
	bge 大于等于时分支, B-Type, RV32I and RV64I, if(x[rs1] >= x[rs2])	pc += sext(imm);
	若寄存器x[rs1]的值大于等于寄存器x[rs2]的值(均视有有符号数)，把pc的值设置为当前值加上符号位扩展的立即数;
	+----------------------------------------------------------------------------+
	|31				 25|24		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|	imm[12|10:5]   |    rs2	  |    rs1    |  101  | imm[4:1|11] |   1100011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_bge = opcode_is_1100011 & funct3_is_101;

/*
	bgeu 无符号大于等于时分支, B-Type, RV32I and RV64I, if(x[rs1] >= x[rs2])	pc += sext(imm);
	若寄存器x[rs1]的值大于等于寄存器x[rs2]的值(均视为无符号数)，把pc的值设置为当前值加上符号位扩展的立即数;
	+----------------------------------------------------------------------------+
	|31				 25|24		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|	imm[12|10:5]   |    rs2	  |    rs1    |  111  | imm[4:1|11] |   1100011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_bgeu = opcode_is_1100011 & funct3_is_111;

/*
	blt 小于时分支，B-Type，RV32I and RV64I，if(x[rs1] < x[rs2])  pc += sext(imm)
	若寄存器x[rs1]的值小于寄存器x[rs2]的值，有符号数，则把pc的值设为当前值加上符号位扩展的立即数;
	+----------------------------------------------------------------------------+
	|31				 25|24		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|	imm[12|10:5]   |    rs2	  |    rs1    |  100  | imm[4:1|11] |   1100011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_blt = opcode_is_1100011 & funct3_is_100;

/*
	bltu 小于时分支，B-Type，RV32I and RV64I，if(x[rs1] < x[rs2])  pc += sext(imm)
	若寄存器x[rs1]的值小于寄存器x[rs2]的值，无符号数，则把pc的值设为当前值加上符号位扩展的立即数;
	+----------------------------------------------------------------------------+
	|31				 25|24		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|	imm[12|10:5]   |    rs2	  |    rs1    |  110  | imm[4:1|11] |   1100011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_bltu = opcode_is_1100011 & funct3_is_110;

/*
	bne 不相等时分支，B-Type，RV32I and RV64I，if(x[rs1] != x[rs2])  pc += sext(imm)
	若寄存器x[rs1]的值不等于寄存器x[rs2]的值，则把pc的值设为当前值加上符号位扩展的立即数;
	+----------------------------------------------------------------------------+
	|31				 25|24		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|	imm[12|10:5]   |    rs2	  |    rs1    |  001  | imm[4:1|11] |   1100011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_bne = opcode_is_1100011 & funct3_is_001;

/*
	csrrc 读后清除控制状态寄存器， t = CSRs[csr]; CSRs[csr] = t & (~x[rs1]); x[rd] = t
	记控制状态寄存器csr中的值为t，把t和寄存器x[rs1]按位与的结果写入csr，两把t写入x[rd]
	+----------------------------------------------------------------------------+
	|31				 			20|19		15|14	12|11		   7|6			0|
	+-----------------------------+-----------+-------+-------------+------------+
	|			csr				  |    rs1    |  011  | 	rd		|   1110011  |
	+----------------------------------------------------------------------------+	
*/
assign      instr_is_csrrc = opcode_is_1110011 & funct3_is_011;

/*
	csrrci 立即数读后清除控制状态寄存器， t = CSRs[csr]; CSRs[csr] = t & (~zimm); x[rd] = t
	记控制状态寄存器csr中的值为t，把t和和五位零扩展的立即数zimm拉位与的结果写入csr，再把t
	写入x[rd](csr寄存器的第五位及更高位不娈)
	+----------------------------------------------------------------------------+
	|31				 			20|19		15|14	12|11		   7|6			0|
	+-----------------------------+-----------+-------+-------------+------------+
	|			csr				  |	zimm[4:0] |  111  | 	rd		|   1110011  |
	+----------------------------------------------------------------------------+	
*/
assign      instr_is_csrrci = opcode_is_1110011 & funct3_is_111;

/*
	csrrs 读后置位控制状态寄存器， t = CSRs[csr]; CSRs[csr] = t | x[rs1]; x[rd] = t
	记控制状态寄存器csr中的值为t，把t和寄存器x[rs1]按位或的结果写入csr，两把t写入x[rd]
	+----------------------------------------------------------------------------+
	|31				 			20|19		15|14	12|11		   7|6			0|
	+-----------------------------+-----------+-------+-------------+------------+
	|			csr				  |    rs1    |  010  | 	rd		|   1110011  |
	+----------------------------------------------------------------------------+	
*/
assign      instr_is_csrrs = opcode_is_1110011 & funct3_is_010;

/*
	csrrsi 立即数读设置控制状态寄存器， t = CSRs[csr]; CSRs[csr] = t | zimm; x[rd] = t
	记控制状态寄存器csr中的值为t，把t和和五位零扩展的立即数zimm拉位或的结果写入csr，再把t
	写入x[rd](csr寄存器的第五位及更高位不娈)
	+----------------------------------------------------------------------------+
	|31				 			20|19		15|14	12|11		   7|6			0|
	+-----------------------------+-----------+-------+-------------+------------+
	|			csr				  |	zimm[4:0] |  110  | 	rd		|   1110011  |
	+----------------------------------------------------------------------------+	
*/
assign      instr_is_csrrsi = opcode_is_1110011 & funct3_is_110;

/*
	csrrw 读后写控制状态寄存器， t = CSRs[csr]; CSRs[csr] = x[rs1]; x[rd] = t
	记控制状态寄存器csr中的值为t，把寄存器x[rs1]的值写入csr，再把t写入x[rd]
	+----------------------------------------------------------------------------+
	|31				 			20|19		15|14	12|11		   7|6			0|
	+-----------------------------+-----------+-------+-------------+------------+
	|			csr				  |		rs1	  |  001  | 	rd		|   1110011  |
	+----------------------------------------------------------------------------+	
*/
assign      instr_is_csrrw = opcode_is_1110011 & funct3_is_001;

/*
	csrrwi 立即数读后写控制状态寄存器， x[rd] = CSRs[csr];CSRs[csr] = zimm
	把控制状态寄存器csr中的值写入x[rd]，再把五位的零扩展的立即数zimm的值写入csr
	+----------------------------------------------------------------------------+
	|31				 			20|19		15|14	12|11		   7|6			0|
	+-----------------------------+-----------+-------+-------------+------------+
	|			csr				  |	zimm[4:0] |  101  | 	rd		|   1110011  |
	+----------------------------------------------------------------------------+	
*/
assign      instr_is_csrrwi = opcode_is_1110011 & funct3_is_101;

/*
	ebreak 环境断点，通过抛出断点异常的方式请求调试器
	+----------------------------------------------------------------------------+
	|31				 			20|19		15|14	12|11		   7|6			0|
	+-----------------------------+-----------+-------+-------------+------------+
	|		000000000001		  |	 00000	  |  000  | 	00000	|   1110011  |
	+----------------------------------------------------------------------------+	
*/
assign      instr_is_ebreak = (ir[31 : 20] == 12'b0000_0000_0001) & funct3_is_000 & opcode_is_1110011;

/*
	ebreak 环境调用，通过引发环境异常的方式请求调试器
	+----------------------------------------------------------------------------+
	|31				 			20|19		15|14	12|11		   7|6			0|
	+-----------------------------+-----------+-------+-------------+------------+
	|		000000000000		  |	 00000	  |  000  | 	00000	|   1110011  |
	+----------------------------------------------------------------------------+	
*/
assign      instr_is_ecall = (ir[31 : 20] == 12'b0000_0000_0000) & funct3_is_000 & opcode_is_1110011;


/*
	fence 同步内存和IO，在后续指令中的内存和IO访问对外部（例如其他线程）可见之前，使这条指令
	之前的内存及IO访问对外部可见，比特中的第3，2，1，0位分别对应设备输入、设备输出、内存读写。
	例如fence r, rw，将前面读取与后面的读取和写入排序，使用pred=0010和succ=0011进行编号。
	如果省略了参数，则表示fence iorw, iorw，即对所有访存请求进行排序。
	+----------------------------------------------------------------------------+
	|31	 	28|27	 24|23		20|19		15|14	12|11		   7|6			0|
	+---------+--------+----------+-----------+-------+-------------+------------+
	| 	0000  | pred   |    succ  |   00000   |  000  | 	00000	|   0001111  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_fence = opcode_is_0001111 & funct3_is_000;

/*
	fencei 同步指令流 使内存指令区域的读写，对后续指令可见
	+----------------------------------------------------------------------------+
	|31	 						20|19		15|14	12|11		   7|6			0|
	+-----------------------------+-----------+-------+-------------+------------+
	| 			000000000000	  |   00000   |  001  | 	00000	|   0001111  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_fencei = opcode_is_0001111 & funct3_is_001;

/*
	jal 跳转并链接 J-Type RV32I and RV64I	x[rd] = pc + 4; pc += sext(imm)
	把下一条指令的地址(pc+4)，然后把pc设置为当前值加上符号位扩展的imm,rd默认为x1
	+----------------------------------------------------------------------------+
	|31	 											12|11		   7|6			0|
	+-------------------------------------------------+-------------+------------+
	| 				imm[20|10:1|11|19:12] 			  | 	rd		|   1101111  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_jal = opcode_is_1101111;

/*
	jalr 跳转并链接寄存器 I-Type	t = pc + 4; pc = (x[rs1] + sext(imm)) & ~1; x[rd] = t
	把pc设置为x[rs1] + sext(imm)，把计算出来的地址的最低有效位设为0，并将原pc+4写入x[rd],rd默认为x1
	+----------------------------------------------------------------------------+
	|31				 			20|19		15|14	12|11		   7|6			0|
	+-----------------------------+-----------+-------+-------------+------------+
	|			imm[11:0]		  |	 	rs1	  |  010  | 	rd		|   1100111  |
	+----------------------------------------------------------------------------+	
*/
assign      instr_is_jalr = opcode_is_1100111 & funct3_is_000;

/*
	lb 字节加载，I-Type RV32I and RV64I		x[rd] = sext(M[x[rs1] + sext(imm)][7:0])
	从地址x[rs1] + sext(imm)处读取一个字节，经符号位扩展后写入x[rd]
	+----------------------------------------------------------------------------+
	|31				 			20|19		15|14	12|11		   7|6			0|
	+-----------------------------+-----------+-------+-------------+------------+
	|			imm[11:0]		  |	 	rs1	  |  000  | 	rd		|   0000011  |
	+----------------------------------------------------------------------------+	
*/
assign      instr_is_lb = opcode_is_0000011 & funct3_is_000;

/*
	lbu 无符号字节加载，I-Type RV32I and RV64I	x[rd] = M[x[rs1] + sext(imm)][7:0]
	从地址x[rs1] + sext(imm)处读取一个字节，经零扩展后写入x[rd]
	+----------------------------------------------------------------------------+
	|31				 			20|19		15|14	12|11		   7|6			0|
	+-----------------------------+-----------+-------+-------------+------------+
	|			imm[11:0]		  |	 	rs1	  |  100  | 	rd		|   0000011  |
	+----------------------------------------------------------------------------+	
*/
assign      instr_is_lbu = opcode_is_0000011 & funct3_is_100;

/*
	lh 半字加载，I-Type RV32I and RV64I	x[rd] = sext(M[x[rs1] + sext(imm)][15:0])
	从地址x[rs1] + sext(imm)处读取两个字节，经符号位扩展后写入x[rd]
	+----------------------------------------------------------------------------+
	|31				 			20|19		15|14	12|11		   7|6			0|
	+-----------------------------+-----------+-------+-------------+------------+
	|			imm[11:0]		  |	 	rs1	  |  001  | 	rd		|   0000011  |
	+----------------------------------------------------------------------------+	
*/
assign      instr_is_lh = opcode_is_0000011 & funct3_is_001;

/*
	lhu 半字加载，I-Type RV32I and RV64I	x[rd] = M[x[rs1] + sext(imm)][15:0]
	从地址x[rs1] + sext(imm)处读取两个字节，经零扩展后写入x[rd]
	+----------------------------------------------------------------------------+
	|31				 			20|19		15|14	12|11		   7|6			0|
	+-----------------------------+-----------+-------+-------------+------------+
	|			imm[11:0]		  |	 	rs1	  |  101  | 	rd		|   0000011  |
	+----------------------------------------------------------------------------+	
*/
assign      instr_is_lhu = opcode_is_0000011 & funct3_is_101;

/*
	lw 字加载，I-Type，RV32I and RV64I，x[rd] = sext(Mem[x[rs1] + sext(imm[11 : 0])][31 : 0]);
	从地址x[rs1] + sign-extend(imm[11 : 0])读取四个字节，写入x[rd]
	+----------------------------------------------------------------------------+
	|31				 			20|19		15|14	12|11		   7|6			0|
	+-----------------------------+-----------+-------+-------------+------------+
	|			imm[11:0]		  |	 	rs1	  |  010  | 	rd		|   0000011  |
	+----------------------------------------------------------------------------+	
*/
assign      instr_is_lw = opcode_is_0000011 & funct3_is_010;

/* 
    lui 高位立即数加载，U Type，RV32I and RV64I，x[rd] = sext(imm[31 : 12] << 12);
    将符号位扩展的20位立即数imm左移12位，并将低12位置0，写入x[rd]中。
    +----------------------------------------------------------------------------+
    |31                                             12|11          7|6          0|
    +-------------------------------------------------+-------------+------------+
    |                   imm[31：12]                   |     rd      |   0110111  |
    +----------------------------------------------------------------------------+
*/
assign      instr_is_lui = opcode_is_0110111;

/*
    mret 机器模式异常返回	R-Type RV32I and RV64I特权架构
    从机器模式异常处理程序返回，将pc设置为CSRs[mepc]，将特权级设置为CSRs[mstatus].MPP，
    CSRs[msatus].MIE设置为CSRs[mstatus].MPIE，并且将CSRs[mstatus].MPIE设置为1；并且，
    如果支持用户模式，则将CSRs[mstatus].MPP设置为0
    +----------------------------------------------------------------------------+
    |31				 25|24		20|19		15|14	12|11		   7|6			0|
    +------------------+----------+-----------+-------+-------------+------------+
    |		0011000	   |  00010	  |    00000  |  000  | 	00000 	|   1110011  |
    +----------------------------------------------------------------------------+
*/
assign      instr_is_mret = (ir[31 : 20] == 12'b0011_0000_0010) & funct3_is_000 & opcode_is_1110011;


/*
    dret 调试模式返回
*/
assign      instr_is_dret = (ir[31 : 20] == 12'b0111_1011_0010) & funct3_is_000 & opcode_is_1110011;

/*
	or 或, R-Type, RV32I and RV64I, 					x[rd] = x[rs1] | x[rs2];
	将寄存器x[rs1]和寄存器x[rs2]位或的结果写入x[rd]寄存器.
	+----------------------------------------------------------------------------+
	|31				 25|24		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|		0000000	   |    rs2	  |    rs1    |  110  | 	rd		|   0110011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_or = opcode_is_0110011 & funct3_is_110 & funct7_is_0000000;

/*
	ori 立即数或, R-Type, RV32I and RV64I, 					x[rd] = x[rs1] | sext(imm);
	将寄存器x[rs1]和寄存器x[rs2]位或的结果写入x[rd]寄存器.
	+----------------------------------------------------------------------------+
	|31				 25|24		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|	imm[11:0]	   |    rs2	  |    rs1    |  110  | 	rd		|   0010011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_ori = opcode_is_0010011 & funct3_is_110;

/*
	sb	存字节	S-Type	RV32I and RV64I			M[x[rs1]+ sext(imm)] = x[rs2][7:0]
	将x[rs2]的低字节存入内存地址x[rs1] + sext(imm)
	+----------------------------------------------------------------------------+
	|31				 25|24		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|	imm[11:5]	   |    rs2	  |    rs1    |  000  | imm[4:0]	|   0100011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_sb = opcode_is_0100011 & funct3_is_000;

/*
	sh	存半字	S-Type	RV32I and RV64I			M[x[rs1]+ sext(imm)] = x[rs2][15:0]
	将x[rs2]的低半字存入内存地址x[rs1] + sext(imm)
	+----------------------------------------------------------------------------+
	|31				 25|24		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|	imm[11:5]	   |    rs2	  |    rs1    |  001  | imm[4:0]	|   0100011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_sh = opcode_is_0100011 & funct3_is_001;

/*
	sh	存字	S-Type	RV32I and RV64I			M[x[rs1]+ sext(imm)] = x[rs2]
	将x[rs2]存入内存地址x[rs1] + sext(imm)
	+----------------------------------------------------------------------------+
	|31				 25|24		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|	imm[11:5]	   |    rs2	  |    rs1    |  010  | imm[4:0]	|   0100011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_sw = opcode_is_0100011 & funct3_is_010;

/*
	sll	逻辑左移 R-Type RV32I and RV64I			x[rd] = x[rs1] << x[rs2]
	把寄存器x[rs1]左移x[rs2]位，空出的位置补0，结果写入x[rd]。x[rs2]的低5位代表移动位数，
	高位忽略
	+----------------------------------------------------------------------------+
	|31				 25|24		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|		0000000	   |    rs2	  |    rs1    |  001  | 	rd		|   0110011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_sll = opcode_is_0110011 & funct3_is_001 & funct7_is_0000000;

/*
	slli	立即数逻辑左移 R-Type RV32I and RV64I			x[rd] = x[rs1] << imm
	把寄存器x[rs1]左移imm位，空出的位置补0，结果写入x[rd]。对于RV32I，仅当imm[5]=0时，
	指令才有效
	+----------------------------------------------------------------------------+
	|31				 26|25		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|		000000	   |    imm	  |    rs1    |  001  | 	rd		|   0010011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_slli = opcode_is_0010011 & funct3_is_001 & funct7_is_0000000;

/*
	slt	小于则置位	R-Type	RV32I and RV64I			x[rd] = x[rs1] < x[rs2]
	比较x[rs1]和x[rs2]中的数，如果x[rs1]更小，向x[rd]写入1，否则写入0
	+----------------------------------------------------------------------------+
	|31				 25|24		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|		0000000	   |    rs2	  |    rs1    |  010  | 	rd		|   0110011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_slt = opcode_is_0110011 & funct3_is_010 & funct7_is_0000000;

/*
	slti 小于立即数则置位	I-Type RV32I and RV64I	x[rd] = x[rs1] < sext(imm)
	比较x[rs1]和有符号扩展的立即数，如果x[rs1]更小，向x[rd]写入1，否则写入0
	+----------------------------------------------------------------------------+
	|31				 			20|19		15|14	12|11		   7|6			0|
	+-----------------------------+-----------+-------+-------------+------------+
	|			imm[11:0]		  |	 	rs1	  |  010  | 	rd		|   0010011  |
	+----------------------------------------------------------------------------+	
*/
assign      instr_is_slti = opcode_is_0010011 & funct3_is_010;

/*
	sltiu 无符号小于立即数则置位	I-Type RV32I and RV64I	x[rd] = x[rs1] < ext(imm)
	比较x[rs1]和零扩展的立即数，比较时视为无符号数，如果x[rs1]更小，向x[rd]写入1，否则
	写入0
	+----------------------------------------------------------------------------+
	|31				 			20|19		15|14	12|11		   7|6			0|
	+-----------------------------+-----------+-------+-------------+------------+
	|			imm[11:0]		  |	 	rs1	  |  011  | 	rd		|   0010011  |
	+----------------------------------------------------------------------------+	
*/
assign      instr_is_sltiu = opcode_is_0010011 & funct3_is_011;

/*
	sltu 无符号小于则置位	R-Type	RV32I and RV64I			x[rd] = x[rs1] < x[rs2]
	比较x[rs1]和x[rs2]中的数，比较时视为无符号数，如果x[rs1]更小，向x[rd]写入1，否则写入0
	+----------------------------------------------------------------------------+
	|31				 25|24		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|		0000000	   |    rs2	  |    rs1    |  011  | 	rd		|   0110011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_sltu = opcode_is_0110011 & funct3_is_011 & funct7_is_0000000;

/*
	sra	算术右移 R-Type RV32I and RV64I			x[rd] = x[rs1] >> x[rs2]
	把寄存器x[rs1]右移x[rs2]位，空位用x[rs1]的最高位填充，结果写入x[rd]。x[rs2]的低5位
	代表移动位数，高位忽略
	+----------------------------------------------------------------------------+
	|31				 25|24		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|		0100000	   |    rs2	  |    rs1    |  101  | 	rd		|   0110011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_sra = opcode_is_0110011 & funct3_is_101 & funct7_is_0100000;

/*
	srai 立即数算术右移 R-Type RV32I and RV64I			x[rd] = x[rs1] >> x[rs2]
	把寄存器x[rs1]右移imm位，空位用x[rs1]的最高位填充，结果写入x[rd]。仅当imm[5]=0时有效
	+----------------------------------------------------------------------------+
	|31				 26|25		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|		010000	   |    imm	  |    rs1    |  101  | 	rd		|   0010011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_srai = opcode_is_0010011 & funct3_is_101 & funct7_is_0100000;

/*
	srl	逻辑右移 R-Type RV32I and RV64I			x[rd] = x[rs1] >> x[rs2]
	把寄存器x[rs1]右移x[rs2]位，空位用0填充，结果写入x[rd]。x[rs2]的低5位代表移动位数，
	高位忽略
	+----------------------------------------------------------------------------+
	|31				 25|24		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|		0000000	   |    rs2	  |    rs1    |  101  | 	rd		|   0110011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_srl = opcode_is_0110011 & funct3_is_101 & funct7_is_0000000;

/*
	srai 立即数逻辑右移 R-Type RV32I and RV64I			x[rd] = x[rs1] >> imm
	把寄存器x[rs1]右移imm位，空位用0填充，结果写入x[rd]。仅当imm[5]=0时有效
	+----------------------------------------------------------------------------+
	|31				 26|25		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|		000000	   |    imm	  |    rs1    |  101  | 	rd		|   0010011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_srli = opcode_is_0010011 & funct3_is_101 & funct7_is_0000000;

/*
	sub 减，R-Type，RV32I and RV64I，	x[rd] = x[rs1] - x[rs2]，忽略算术溢出
	+----------------------------------------------------------------------------+
	|31				 25|24		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|		0100000	   |    rs2	  |    rs1    |  000  | 	rd		|   0110011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_sub = opcode_is_0110011 & funct3_is_000 & funct7_is_0100000;

/*
	wfi 特权指令，等待中断，如果没有待处理的中断，则将处理器置为空闲状态
	+----------------------------------------------------------------------------+
	|31				 25|24		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|		0001000	   |   00101  |   00000   |  000  | 	00000	|   1110011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_wfi = funct7_is_0001000 & funct3_is_000 & opcode_is_1110011;

/*
	xor 异或, R-Type, RV32I and RV64I, 					x[rd] = x[rs1] ^ x[rs2];
	将寄存器x[rs1]和寄存器x[rs2]异或的结果写入x[rd]寄存器.
	+----------------------------------------------------------------------------+
	|31				 25|24		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|		0000000	   |    rs2	  |    rs1    |  100  | 	rd		|   0110011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_xor = opcode_is_0110011 & funct3_is_100 & funct7_is_0000000;

/*
	xori 立即数异或, R-Type, RV32I and RV64I, 			x[rd] = x[rs1] ^ sext(imm);
	将寄存器x[rs1]和寄存器x[rs2]异或的结果写入x[rd]寄存器.
	+----------------------------------------------------------------------------+
	|31				 25|24		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|	imm[11:0]	   |    rs2	  |    rs1    |  100  | 	rd		|   0010011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_xori = opcode_is_0010011 & funct3_is_100;


/*
	div 除法 R-Type, Rv32M and RV64M, x[rd] = x[rs1] / x[rs2]；
	用寄存器x[rs1]的值除以寄存器x[rs2]的值，向零舍入，将这些数视为二进制补码，把商写入x[rd]
	+----------------------------------------------------------------------------+
	|31				 25|24		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|		0000001	   |    rs2	  |    rs1    |  100  | 	rd		|   0110011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_div = opcode_is_0110011 & funct3_is_100 & funct7_is_0000001;

/*
	divu 无符号除法 R-Type, Rv32M and RV64M, x[rd] = x[rs1] / x[rs2]；
	用寄存器x[rs1]的值除以寄存器x[rs2]的值，向零舍入，将这些数视为无符号数，把商写入x[rd]
	+----------------------------------------------------------------------------+
	|31				 25|24		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|		0000001	   |    rs2	  |    rs1    |  101  | 	rd		|   0110011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_divu = opcode_is_0110011 & funct3_is_101 & funct7_is_0000001;

/*
	mul	乘 R-Type RV32I and RV64I，						x[rd] = x[rs1] * x[rs2]
	把寄存器x[rs1]与寄存器x[rs2]的乘积写入x[rd]，忽略算术溢出
	+----------------------------------------------------------------------------+
	|31				 25|24		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|		0000001	   |    rs2	  |    rs1    |  000  | 	rd		|   0110011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_mul = opcode_is_0110011 & funct3_is_000 & funct7_is_0000001;

/*
	mulh 高位乘 R-Type RV32I and RV64I，			x[rd] = x[rs1] * x[rs2] >> XLEN
	将寄存器x[rs1]与寄存器x[rs2]相乘，x[rs1]、x[rs2]都视为二进制补码，将乘积的高位写入x[rd]
	+----------------------------------------------------------------------------+
	|31				 25|24		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|		0000001	   |    rs2	  |    rs1    |  001  | 	rd		|   0110011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_mulh = opcode_is_0110011 & funct3_is_001 & funct7_is_0000001;

/*
	mulhsu 高位乘 R-Type RV32I and RV64I，			x[rd] = x[rs1] * x[rs2] >> XLEN
	将寄存器x[rs1]与寄存器x[rs2]相乘，x[rs1]为二进制补码，x[rs2]为无符号数，将乘积的高位
	写入x[rd]
	+----------------------------------------------------------------------------+
	|31				 25|24		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|		0000001	   |    rs2	  |    rs1    |  010  | 	rd		|   0110011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_mulhsu = opcode_is_0110011 & funct3_is_010 & funct7_is_0000001;

/*
	mulhu 高位无符号乘 R-Type RV32I and RV64I，			x[rd] = x[rs1] * x[rs2] >> XLEN
	将寄存器x[rs1]与寄存器x[rs2]相乘，x[rs1]、x[rs2]都视为无符号数，将乘积的高位写入x[rd]
	+----------------------------------------------------------------------------+
	|31				 25|24		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|		0000001	   |    rs2	  |    rs1    |  001  | 	rd		|   0110011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_mulhu = opcode_is_0110011 & funct3_is_011 & funct7_is_0000001;

/*
	rem	求余数 R-Type RV32I and RV64I，						x[rd] = x[rs1] % x[rs2]
	x[rs1]除以x[rs2]，向0舍入，都视为二进制数，余数写入x[rd]
	+----------------------------------------------------------------------------+
	|31				 25|24		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|		0000001	   |    rs2	  |    rs1    |  110  | 	rd		|   0110011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_rem = opcode_is_0110011 & funct3_is_110 & funct7_is_0000001;

/*
	rem	求无符号的余数 R-Type RV32I and RV64I，				x[rd] = x[rs1] % x[rs2]
	x[rs1]除以x[rs2]，向0舍入，都视为无符号数，余数写入x[rd]
	+----------------------------------------------------------------------------+
	|31				 25|24		20|19		15|14	12|11		   7|6			0|
	+------------------+----------+-----------+-------+-------------+------------+
	|		0000001	   |    rs2	  |    rs1    |  111  | 	rd		|   0110011  |
	+----------------------------------------------------------------------------+
*/
assign      instr_is_remu = opcode_is_0110011 & funct3_is_111 & funct7_is_0000001;



/*********************************** 指令立即数解析/选择部分 ****************************************/
/*
	对于U型指令，需要操作立即数的指令：lui auipc
	J型指令，只有jal指令需要操作立即数;
	B型指令都需要操作立即数;
	I型指令部分需要操作立即数，其中slli、srli、srali的立即数与其他指令的位置不一样，需要单独处理;
	S型
*/
// 从指令中解析出立即数
assign      i_type_imm      = `GET_I_TYPE_IMM(ir);
assign      i_type_shamt    = `GET_I_TYPE_SHAMT(ir);
assign      i_type_zimm     = `GET_I_TYPE_ZIMM(ir);
assign      b_type_bxx_imm  = `GET_B_TYPE_BXX_IMM(ir);
assign      b_type_jal_imm  = `GET_B_TYPE_JAL_IMM(ir);
assign      s_type_imm      = `GET_S_TYPE_IMM(ir);
assign      u_type_imm      = `GET_U_TYPE_IMM(ir);

assign      sel_i_type_imm =    opcode_is_0010011  | 
                                instr_is_jalr | 
                                opcode_is_0000011;

// csrrci csrrsi csrrwi需要使用zimm
assign      sel_i_type_zimm = opcode_is_1110011 & 
                                (
                                    funct3_is_101 | 
                                    funct3_is_110 | 
                                    funct3_is_111
                                );

assign      sel_b_type_bxx_imm = opcode_is_1100011;

assign      sel_b_type_jal_imm = instr_is_jal;

assign      sel_s_type_imm = opcode_is_0100011;

assign      sel_u_type_imm = instr_is_lui | instr_is_auipc;


// 选择立即数输出
assign      dec_imm =   ({32{sel_i_type_imm     }} & i_type_imm         ) | 
                        ({32{sel_i_type_zimm    }} & i_type_zimm        ) | 
                        ({32{sel_b_type_bxx_imm }} & b_type_bxx_imm     ) | 
                        ({32{sel_b_type_jal_imm }} & b_type_jal_imm     ) | 
                        ({32{sel_s_type_imm     }} & s_type_imm         ) | 
                        ({32{sel_u_type_imm     }} & u_type_imm         );



// 将指令分为以下几类
// 1、常规运算指令，包含:
//      add addi auipc sub and andi or ori xor xori lui sll slli slt slti sltu sltiu sra srai srl srli
// 2、分支指令，包含:
//      beq bge bgeu blt bltu bne jal jalr mret dret
// 3、系统相关指令，包含:
//      ebreak ecall fence fencei wfi csrrc csrrci csrrw csrrwi csrrs csrrsi
// 4、lsu指令，需要访存，包含:
//      lb lbu lh lhu lw sb sh sw
// 5、乘除法指令，包含:
//      div divu mul mulh mulhsu mulhu rem remu
// 6、原子指令，需要访存
//
// 7、浮点运算指令

// 常规运算指令
assign      rglr_op_bus[`RGLR_ADD_LOC]      = instr_is_add | instr_is_addi;
assign      rglr_op_bus[`RGLR_SUB_LOC]      = instr_is_sub;
assign      rglr_op_bus[`RGLR_AND_LOC]      = instr_is_and | instr_is_andi;
assign      rglr_op_bus[`RGLR_OR_LOC]       = instr_is_or | instr_is_ori;
assign      rglr_op_bus[`RGLR_XOR_LOC]      = instr_is_xor | instr_is_xori;
assign      rglr_op_bus[`RGLR_SLL_LOC]      = instr_is_sll | instr_is_slli;
assign      rglr_op_bus[`RGLR_SLT_LOC]      = instr_is_slt | instr_is_slti;
assign      rglr_op_bus[`RGLR_SRA_LOC]      = instr_is_sra | instr_is_srai;
assign      rglr_op_bus[`RGLR_SRL_LOC]      = instr_is_srl | instr_is_srli;
assign      rglr_op_bus[`RGLR_AUIPC_LOC]    = instr_is_auipc;
assign      rglr_op_bus[`RGLR_LUI_LOC]      = instr_is_lui;
assign      rglr_op_bus[`RGLR_SLTU_LOC]     = instr_is_sltu | instr_is_sltiu;
assign      rglr_op_bus[`RGLR_OP1_IS_PC]    = instr_is_auipc;
assign      rglr_op_bus[`RGLR_OP2_IS_IMM]   = instr_is_i_type | instr_is_u_type;
assign      dec_rglr_instr =    opcode_is_0010011 | 
                                (opcode_is_0110011 & (~funct7_is_0000001)) | 	//opcode == 0110011 且 funct7 == 0000001时，为乘除法指令
                                instr_is_lui | 
                                instr_is_auipc;


// 访存指令
assign      lsu_op_bus[`LSU_LOAD_LOC]   = instr_is_lb | instr_is_lh | instr_is_lw | instr_is_lbu | instr_is_lhu;
assign      lsu_op_bus[`LSU_STORE_LOC]  = instr_is_sb | instr_is_sh | instr_is_sw;
assign      lsu_op_bus[`LSU_SIZE_LOC]   =   (instr_is_lb | instr_is_lbu | instr_is_sb) ?  2'd0 : 
                                            (instr_is_lh | instr_is_lhu | instr_is_sh) ? 2'd1 : 
                                            2'd2;
assign      lsu_op_bus[`LSU_UEXT_LOC]   = instr_is_lbu | instr_is_lhu;
assign      dec_lsu_instr = opcode_is_0000011 | 
                            opcode_is_0100011 | 
`ifdef  LNRV_SUPPORTED_AMO
                            opcode_is_0101111 | 
`endif
                            1'b0;


// 分支指令
assign      brch_op_bus[`BRCH_BEQ_LOC]      = instr_is_beq;
assign      brch_op_bus[`BRCH_BGE_LOC]      = instr_is_bge;
assign      brch_op_bus[`BRCH_BGEU_LOC]     = instr_is_bgeu;
assign      brch_op_bus[`BRCH_BLT_LOC]      = instr_is_blt;
assign      brch_op_bus[`BRCH_BLTU_LOC]     = instr_is_bltu;
assign      brch_op_bus[`BRCH_BNE_LOC]      = instr_is_bne;
assign      brch_op_bus[`BRCH_JAL_LOC]      = instr_is_jal;
assign      brch_op_bus[`BRCH_JALR_LOC]     = instr_is_jalr;
assign      brch_op_bus[`BRCH_MRET_LOC]     = instr_is_mret;
assign      brch_op_bus[`BRCH_DRET_LOC]     = instr_is_dret;
assign      brch_op_bus[`BRCH_FENCE_LOC]    = instr_is_fence | instr_is_fencei;
assign      brch_op_bus[`BRCH_OP1_IS_PC]    = instr_is_jal | instr_is_jalr;
assign      brch_op_bus[`BRCH_OP2_IS_IMM] = instr_is_jal | instr_is_jalr;
assign      dec_brch_instr  = opcode_is_1100011 | 
                                instr_is_jal |
                                instr_is_jalr | 
                                instr_is_mret | 
                                legl_dret;


// csr操作指令
assign      csr_op_bus[`CSR_CSRRC_LOC] = instr_is_csrrc | instr_is_csrrci;
assign      csr_op_bus[`CSR_CSRRS_LOC] = instr_is_csrrs | instr_is_csrrsi;
assign      csr_op_bus[`CSR_CSRRW_LOC] = instr_is_csrrw | instr_is_csrrwi;
assign      csr_op_bus[`CSR_OP1_IS_ZERO] = csr_op_bus[`CSR_CSRRS_LOC];
assign      csr_op_bus[`CSR_OP2_IS_IMM] = instr_is_csrrci | instr_is_csrrsi | instr_is_csrrwi;
assign      dec_csr_instr = opcode_is_1110011 & (~funct3_is_000);

// 系统相关指令
assign      sys_op_bus[`SYS_WFI_LOC] = instr_is_wfi;
assign      sys_op_bus[`SYS_EBREAK_LOC] = instr_is_ebreak;
assign      sys_op_bus[`SYS_ECALL_LOC] = instr_is_ecall;
assign      dec_sys_instr = instr_is_wfi | 
                            instr_is_ebreak | 
                            instr_is_ecall;


/* 如果存在乘法/除法单元则需要译码相关指令 */

// 乘法相关指令
assign      mdv_op_bus[`MDV_DIV_LOC] = instr_is_div | instr_is_divu;
assign      mdv_op_bus[`MDV_MUL_LOC] = instr_is_mul | instr_is_mulh | instr_is_mulhsu | instr_is_mulhu;
assign      mdv_op_bus[`MDV_REM_LOC] = instr_is_rem | instr_is_remu;
assign      mdv_op_bus[`MDV_OP1_UNSIGNED_LOC] = instr_is_divu | instr_is_mulhu | instr_is_remu;
assign      mdv_op_bus[`MDV_OP2_UNSIGNED_LOC] = instr_is_divu | instr_is_mulhsu | instr_is_mulhu | instr_is_remu;
assign      mdv_op_bus[`MDV_RES_HIGH_LOC] = instr_is_mulh | instr_is_mulhsu | instr_is_mulhu;
assign      dec_mdv_instr = opcode_is_0110011 & funct7_is_0000001;


// 暂时不支持原子指令
assign      dec_amo_instr = 1'b0;

// 暂时不支持浮点运算指令
assign      dec_fpu_instr = 1'b0;

// 选出一个译码信息，由于OP_BUS_WIDTH使用的是各个OP_BUS_WIDTH中最大的那个，如果直接使用OP_BUS_WIDTH - RGLR_OP_BUS_WIDTH，
// 有可能出现{0{1'b0}}的情况，为了避免这个情况发生，我们将op_bus_mux的位宽定义为OP_BUS_WIDTH+1，这样可以保证相减后至少为1,
// 只需要在输出的时候忽略最高位即可。
assign      dec_op_bus_mux =    ({(`DEC_OP_BUS_WIDTH + 1){dec_rglr_instr}} & {{(`DEC_OP_BUS_WIDTH + 1 - `RGLR_OP_BUS_WIDTH){1'b0}}, rglr_op_bus}) | 
                                ({(`DEC_OP_BUS_WIDTH + 1){dec_brch_instr}} & {{(`DEC_OP_BUS_WIDTH + 1 - `BRCH_OP_BUS_WIDTH){1'b0}}, brch_op_bus}) | 
                                ({(`DEC_OP_BUS_WIDTH + 1){dec_lsu_instr}} & {{(`DEC_OP_BUS_WIDTH + 1 - `LSU_OP_BUS_WIDTH){1'b0}}, lsu_op_bus}) | 
                                ({(`DEC_OP_BUS_WIDTH + 1){dec_csr_instr}} & {{(`DEC_OP_BUS_WIDTH + 1 - `CSR_OP_BUS_WIDTH){1'b0}}, csr_op_bus}) | 
                                ({(`DEC_OP_BUS_WIDTH + 1){dec_sys_instr}} & {{(`DEC_OP_BUS_WIDTH + 1 - `SYS_OP_BUS_WIDTH){1'b0}}, sys_op_bus}) | 
                                ({(`DEC_OP_BUS_WIDTH + 1){dec_mdv_instr}} & {{(`DEC_OP_BUS_WIDTH + 1 - `MDV_OP_BUS_WIDTH){1'b0}}, mdv_op_bus});

assign      dec_op_bus = dec_op_bus_mux[0 +: `DEC_OP_BUS_WIDTH];

// 判断非法指令

// shamt只有在比特5为0的情况下才有效
assign      ilegl_shamt = i_type_shamt[5];
// 
assign      ilegl_sxxi = ilegl_shamt & (instr_is_srai | instr_is_srli | instr_is_slli);

// dret指令只在debug mode下才可以使用
assign      ilegl_dret = instr_is_dret & (~d_mode);
assign      legl_dret = instr_is_dret & d_mode;

// 如果找不到执行模块，也认为是非法指令
assign      legl_exu =  dec_rglr_instr | 
                        dec_sys_instr | 
                        dec_brch_instr | 
                        dec_lsu_instr | 
                        dec_mdv_instr | 
                        dec_fpu_instr | 
                        dec_csr_instr |
                        dec_amo_instr;

assign      ilegl_exu = ~legl_exu;

assign      dec_ilegl_instr =   ilegl_exu |
                                ilegl_sxxi | 
                                ilegl_dret;


assign      dec_rs1_idx = rs1_idx;
assign      dec_rs2_idx = rs2_idx;
assign      dec_rd_idx = rd_idx;
assign      dec_csr_idx = csr_idx;

assign      dec_rv32 = 1'b1;
assign      dec_rv16 = 1'b0;

endmodule