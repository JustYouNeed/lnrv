module lnrv_core_tb;



endmodule