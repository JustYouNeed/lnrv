module lnrv_icb2axi#
(
    parameter                   P_ADDR_WIDTH = 32,
    parameter                   P_DATA_WIDTH = 32
)
(
    input                       clk
);


endmodule