module lnrv_ifu_tb;


endmodule